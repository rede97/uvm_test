module example(input clk);

endmodule